module top(_01_, _07_, _10_, clk, _53_, _73_, _75_, _77_, _79_, _81_, _83_, _85_, _87_, _89_, _91_);
  input  _01_;
  input  _07_;
  input  _10_;
  input  clk;
  output _53_;
  output _73_;
  output _75_;
  output _77_;
  output _79_;
  output _81_;
  output _83_;
  output _85_;
  output _87_;
  output _89_;
  output _91_;
  wire   _03_;
  wire   _09_;
  wire   _13_;
  wire   _18_;
  wire   _20_;
  wire   _21_;
  wire   _22_;
  wire   _24_;
  wire   _25_;
  wire   _33_;
  wire   _62_;
  wire   _63_;
  wire   _64_;
  wire   _65_;
  wire   _66_;
  wire   _67_;
  wire   _68_;
  wire   _69_;
  wire   _70_;
  wire   _71_;
  IBUF _02_ (
    .I(_01_),
    .O(_03_)
  );
  IBUF _08_ (
    .I(_07_),
    .O(_09_)
  );
  IBUF _12_ (
    .I(_10_),
    .O(_13_)
  );
  CARRY4 _16_ (
    .CI(_09_),
    .CYINIT(_09_),
    .DI({_13_, _09_, _03_, _09_}),
    .S({_03_, _03_, _13_, _13_}),
    .CO({_62_, _18_, _63_, _20_}),
    .O({_21_, _22_, _64_, _24_})
  );
  MUXF5 _26_ (
    .I0(_24_),
    .I1(_18_),
    .S(_22_),
    .O(_25_)
  );
  CARRY4 _29_ (
    .CI(_22_),
    .CYINIT(_13_),
    .DI({_21_, _24_, _25_, _22_}),
    .S({_20_, _22_, _09_, _25_}),
    .CO({_65_, _66_, _67_, _33_}),
    .O({_68_, _69_, _70_, _71_})
  );
  OBUF _52_ (
    .I(_33_),
    .O(_53_)
  );
  OBUF _72_ (
    .I(_62_),
    .O(_73_)
  );
  OBUF _74_ (
    .I(_63_),
    .O(_75_)
  );
  OBUF _76_ (
    .I(_64_),
    .O(_77_)
  );
  OBUF _78_ (
    .I(_65_),
    .O(_79_)
  );
  OBUF _80_ (
    .I(_66_),
    .O(_81_)
  );
  OBUF _82_ (
    .I(_67_),
    .O(_83_)
  );
  OBUF _84_ (
    .I(_68_),
    .O(_85_)
  );
  OBUF _86_ (
    .I(_69_),
    .O(_87_)
  );
  OBUF _88_ (
    .I(_70_),
    .O(_89_)
  );
  OBUF _90_ (
    .I(_71_),
    .O(_91_)
  );
endmodule
