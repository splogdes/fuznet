module top(_04_, clk, _12_, _31_, _48_, _50_, _52_, _54_, _56_, _58_, _60_);
  input  _04_;
  input  clk;
  input  _12_;
  output _31_;
  output _48_;
  output _50_;
  output _52_;
  output _54_;
  output _56_;
  output _58_;
  output _60_;
  wire   _03_;
  wire   _07_;
  wire   _11_;
  wire   _14_;
  wire   _19_;
  wire   _40_;
  wire   _41_;
  wire   _42_;
  wire   _43_;
  wire   _44_;
  wire   _45_;
  wire   _46_;
  IBUF _06_ (
    .I(_04_),
    .O(_07_)
  );
  IBUF _13_ (
    .I(_12_),
    .O(_14_)
  );
  CARRY4 _15_ (
    .CI(1'b1),
    .CYINIT(_14_),
    .DI({_07_, _07_, _07_, _14_}),
    .S({_07_, _07_, _07_, _07_}),
    .CO({_40_, _41_, _42_, _19_}),
    .O({_43_, _44_, _45_, _46_})
  );
  OBUF _30_ (
    .I(_19_),
    .O(_31_)
  );
  OBUF _47_ (
    .I(_40_),
    .O(_48_)
  );
  OBUF _49_ (
    .I(_41_),
    .O(_50_)
  );
  OBUF _51_ (
    .I(_42_),
    .O(_52_)
  );
  OBUF _53_ (
    .I(_43_),
    .O(_54_)
  );
  OBUF _55_ (
    .I(_44_),
    .O(_56_)
  );
  OBUF _57_ (
    .I(_45_),
    .O(_58_)
  );
  OBUF _59_ (
    .I(_46_),
    .O(_60_)
  );
endmodule
