module top(_04_, clk, _12_, _31_, _48_, _50_, _52_, _54_, _56_, _58_, _60_);
  input  _04_, _12_;
  input  clk;

  output _31_, _48_, _50_, _52_;
  output _54_, _56_, _58_, _60_;

  wire   _07_, _14_, _19_, _40_, _41_;
  wire   _42_, _43_, _44_, _45_, _46_;

  IBUF _06_ (
    .I(_04_),
    .O(_07_)
  );

  IBUF _13_ (
    .I(_12_),
    .O(_14_)
  );

  CARRY4 _15_ (
    .CI(1'b1),
    .CYINIT(_14_),
    .DI({_07_, _07_, _07_, _14_}),
    .S({_07_, _07_, _07_, _07_}),
    .CO({_40_, _41_, _42_, _19_}),
    .O({_43_, _44_, _45_, _46_})
  );

  OBUF _30_ (
    .I(_19_),
    .O(_31_)
  );

  OBUF _47_ (
    .I(_40_),
    .O(_48_)
  );

  OBUF _49_ (
    .I(_41_),
    .O(_50_)
  );

  OBUF _51_ (
    .I(_42_),
    .O(_52_)
  );

  OBUF _53_ (
    .I(_43_),
    .O(_54_)
  );

  OBUF _55_ (
    .I(_44_),
    .O(_56_)
  );

  OBUF _57_ (
    .I(_45_),
    .O(_58_)
  );

  OBUF _59_ (
    .I(_46_),
    .O(_60_)
  );

endmodule
