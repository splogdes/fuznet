module top(
  input  _005_,
  input  _011_,
  input  _014_,
  input  _015_,
  input  _999_,
  input  clk,
  output _091_,
  output _097_,
  output _101_
);

  wire _003_, _007_, _013_, _017_, _019_, _029_;
  wire _061_, _062_, _064_, _066_, _067_;

  IBUF _006_ (
    .I(_005_),
    .O(_007_)
  );

  IBUF _012_ (
    .I(_011_),
    .O(_013_)
  );

  IBUF _016_ (
    .I(_014_),
    .O(_017_)
  );

  IBUF _072_ (
    .I(_015_),
    .O(_003_)
  );

  IBUF _071_ (
    .I(_999_),
    .O(_029_)
  );

  BUFG _018_ (
    .I(clk),
    .O(_019_)
  );

  SRLC16 #(
    .INIT(16'b0110011001010101)
  ) _060_ (
    .A0(_017_),
    .A1(_017_),
    .A2(_013_),
    .A3(_013_),
    .CLK(_019_),
    .D(_013_),
    .Q(_061_),
    .Q15(_062_)
  );

  LUT1 #(
    .INIT(2'b11)
  ) _898_ (
    .I0(_061_),
    .O(_064_)
  );

  SRLC16 #(
    .INIT(16'b0000011110100000)
  ) _065_ (
    .A0(_003_),
    .A1(_062_),
    .A2(_003_),
    .A3(_007_),
    .CLK(_019_),
    .D(_029_),
    .Q(_066_),
    .Q15(_067_)
  );

  OBUF _090_ (
    .I(_067_),
    .O(_091_)
  );

  OBUF _096_ (
    .I(_066_),
    .O(_097_)
  );

  OBUF _100_ (
    .I(_064_),
    .O(_101_)
  );

endmodule
